module add(input left, input right, output num);
    num = left + right;
endmodule