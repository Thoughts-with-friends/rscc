module add(input a, input b, output num);
    num = a + b;
endmodule
